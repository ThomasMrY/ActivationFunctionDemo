module tanh_1_4_6(x,y);
input wire[5:0]x;
output wire[4:0]y;
assign y[0]=0;
assign y[1]=(x[1]&x[4])|(x[0])|(x[1]&x[3])|(x[1]&x[2]);
assign y[2]=(~x[1]&x[2]&x[5])|(~x[1]&x[2]&x[4])|(~x[1]&x[2]&x[3])|(x[1]&~x[2]&~x[3]&~x[4])|(x[0]);
assign y[3]=(~x[0]&~x[1]&x[3]&x[5])|(~x[0]&~x[1]&x[3]&x[4])|(~x[0]&x[2]&~x[3]&~x[4]&~x[5])|(x[1]&~x[3]&~x[4])|(x[0]&x[1])|(x[1]&x[2])|(x[0]&x[2]&x[3]);
assign y[4]=(~x[0]&~x[1]&x[3]&~x[4]&~x[5])|(~x[0]&x[1]&~x[2]&~x[3]&~x[4])|(~x[0]&x[1]&x[3]&x[4])|(x[0]&~x[1]&~x[2]&x[3]&x[5])|(x[0]&~x[1]&~x[2]&x[3]&x[4])|(x[0]&x[2]&~x[3])|(x[1]&x[2]&x[3])|(~x[2]&x[3]&x[4]&x[5])|(x[2]&~x[3]&x[4]&x[5])|(~x[0]&x[1]&x[3]&x[5])|(~x[0]&~x[1]&~x[2]&x[4]&x[5])|(~x[0]&~x[1]&x[2]&~x[4]&~x[5]);
endmodule