module tanh_1_6_4(x,y);
input wire[3:0]x;
output wire[6:0]y;
assign y[0]=0;
assign y[1]=(x[1]&x[3])|(x[1]&x[2])|(x[0]);
assign y[2]=(~x[1]&x[2]&x[3])|(x[1]&~x[2]&~x[3])|(x[0]);
assign y[3]=(~x[0]&x[2]&~x[3])|(x[1]&~x[3])|(x[1]&x[2])|(x[0]&x[2]&x[3])|(x[0]&x[1]);
assign y[4]=(~x[0]&~x[1]&x[3])|(~x[0]&x[1]&~x[2]&~x[3])|(~x[1]&x[2]&~x[3])|(x[1]&x[2]&x[3])|(x[0]&x[2]&~x[3]);
assign y[5]=(~x[2]&x[3])|(~x[1]&x[2]&~x[3])|(~x[0]&~x[1]&x[3]);
assign y[6]=(~x[2]&x[3])|(~x[0]&~x[1]&x[2]&~x[3])|(x[1]&~x[2])|(x[1]&x[3]);
endmodule